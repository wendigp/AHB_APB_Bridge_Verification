class ahb_agent extends uvm_agent;

	`uvm_component_utils(ahb_agent)

//HANDLE DECLARATIONs
	h_monitor 	monh;
	h_driver	drvh;
	h_sequencer 	seqrh;
	ahb_config	h_cfg;

	extern function new(string name = "ahb_agent", uvm_component parent);
	extern function void build_phase(uvm_phase phase);
	extern function void connect_phase(uvm_phase phase);
endclass

//CONSTRUCTOR
function ahb_agent::new(string name = "ahb_agent", uvm_component parent);
	super.new(name,parent);
endfunction

//BUILD PHASE
function void ahb_agent::build_phase(uvm_phase phase);
	super.build_phase(phase);

	if(!uvm_config_db #(ahb_config)::get(this,"","ahb_config",h_cfg))
	begin
	`uvm_fatal("AHB_AGENT","CANNOT GET DATA FROM AHB_CFG> HAVE YOU SET IT?")
	end

	monh=h_monitor::type_id::create("monh",this);
	
	if(h_cfg.is_active == UVM_ACTIVE)
	begin
	drvh=h_driver::type_id::create("drvh",this);
	seqrh=h_sequencer::type_id::create("seqrh",this);
	end
endfunction

//CONNECT PHASE
function void ahb_agent::connect_phase(uvm_phase phase);
	super.connect_phase(phase);

//CONNECTION OF DRIVER AND SEQUENCER
	if(h_cfg.is_active==UVM_ACTIVE)
	drvh.seq_item_port.connect(seqrh.seq_item_export);
endfunction