class p_monitor extends uvm_monitor;

	`uvm_component_utils(p_monitor)

	virtual apb_if.APB_MON_MP 	vif;
	apb_config 			p_cfg;
	
	uvm_analysis_port#(p_xtn)	monitor_port;

	extern function new(string name = "p_monitor", uvm_component parent);
	extern function void build_phase(uvm_phase phase);
	extern function void connect_phase(uvm_phase phase);
	extern task run_phase(uvm_phase phase);
	extern task collect_data();
endclass

//CONSTRUCTOR
function p_monitor::new(string name = "p_monitor", uvm_component parent);
	super.new(name,parent);
	monitor_port = new("monitor_port",this);
endfunction

//APB MONITOR BUILD PHASE

function void p_monitor::build_phase(uvm_phase phase);
	super.build_phase(phase);

	if(!uvm_config_db #(apb_config)::get(this,"","apb_config",p_cfg))
	begin
	`uvm_fatal("APB MONITOR","CANNOT GET DATA FROM APB_CONFIG. HAVE YOU SET IT?")
	end
endfunction

//APB MONITOR CONNECT PHASE
function void p_monitor::connect_phase(uvm_phase phase);
	super.connect_phase (phase);

	vif = p_cfg.vif;
	if(vif==null)
	begin
	`uvm_fatal("APB_MONITOR","VIF IS NULL IN APB MONITOR")
	end

endfunction

//APB MONITOR RUN PHASE
task p_monitor::run_phase(uvm_phase phase);
	super.run_phase(phase);

	wait(vif.apb_mon_cb.pselx)
	forever
	collect_data();
endtask

task p_monitor::collect_data();

	p_xtn xtn;
	xtn=p_xtn::type_id::create("xtn");

	wait(vif.apb_mon_cb.penable == 1)
	//while(vif.apb_mon_cb.penable != 1)
	//@(vif.apb_mon_cb);
	xtn.paddr = vif.apb_mon_cb.paddr;
	xtn.pwrite = vif.apb_mon_cb.pwrite;
	xtn.penable = vif.apb_mon_cb.penable;
	xtn.pselx = vif.apb_mon_cb.pselx;
	
	if(vif.apb_mon_cb.pwrite == 1)
	xtn.pwdata = vif.apb_mon_cb.pwdata;
	else
	xtn.prdata = vif.apb_mon_cb.prdata;

	`uvm_info("APB MONITOR",$sformatf("Printing from APB MONITOR \n %s",xtn.sprint()), UVM_LOW)
	
	monitor_port.write(xtn);    //SENDS DATA TO SCOREBOARD

	//WAIT FOR TWO CLK CYCLES BEFORE GETTING INTO NEW LOOP - AVOID OVERLAPPING OR GLITCH TRANSACTIONS
	repeat(2) 
	@(vif.apb_mon_cb);
endtask