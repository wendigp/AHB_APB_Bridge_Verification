package test_pkg;



	import uvm_pkg::*;
	`include "uvm_macros.svh"
//	`include "tb_defs.sv"
	`include "h_xtn.sv"
	`include "ahb_config.sv"
	`include "apb_config.sv"
	`include "env_config.sv"
	`include "h_driver.sv"
	`include "h_monitor.sv"
	`include "h_sequencer.sv"
	`include "ahb_agent.sv"
	`include "h_sequence.sv"

	`include "p_xtn.sv"
	`include "p_driver.sv"
	`include "p_monitor.sv"
	`include "p_sequencer.sv"
	`include "apb_agent.sv"
	`include "p_sequence.sv"

	`include "virtual_sequencer.sv"
	`include "virtual_sequence.sv"
	`include "scoreboard.sv"

	`include "env.sv"


	`include "test.sv"
	
endpackage

