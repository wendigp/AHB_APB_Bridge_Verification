class p_xtn extends uvm_sequence_item;

	`uvm_object_utils(p_xtn)

//DECLARATION OF APB PROPERTY
	bit [31:0] paddr;
	bit [31:0] pwdata;
	bit [3:0]  pselx;
	bit		pwrite;
	bit 		penable;
	rand bit [31:0] prdata;

	extern function new(string name = "p_xtn");
	extern function void do_print(uvm_printer printer);

endclass

//CONSTRUCTOR
function p_xtn::new(string name = "p_xtn");
	super.new(name);
endfunction

//PRINT METHOD
function void p_xtn::do_print(uvm_printer printer);
	super.do_print(printer);
	printer.print_field("PADDR",this.paddr,32,UVM_HEX);
	printer.print_field("PWDATA",this.pwdata,32,UVM_HEX);
	printer.print_field("PRDATA",this.prdata,32,UVM_HEX);
	printer.print_field("PSELx",this.pselx,4,UVM_DEC);
	printer.print_field("PWRITE",this.pwrite,1,UVM_BIN);
	printer.print_field("PENABLE",this.penable,1,UVM_BIN);
endfunction